-- this is vga_controller.vhd


















