-- this is top.vhd


