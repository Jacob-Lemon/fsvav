-- this is pixel_generation.vhd

